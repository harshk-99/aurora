module inst_memory (
  input clk,
  input [7:0] mem_address,
  output reg [31:0] data_out
);

integer i;

reg [31:0] rom [256:0];

initial  
      begin                    
                     rom[0]      = 32'b00000000000000000011000000000011;
                     rom[1]      = 32'b00000000000100000011000010000011;
                     rom[2]      = 32'b00000000001000000011000100000011;
                     rom[3]      = 32'b00000000001100000011000110000011;
                     rom[4]      = 32'b00000000010000000011001000000011;
                     rom[5]      = 32'b00000000000000000110000010010011;
                     rom[6]      = 32'b00000000000000000110000100010011;
                     rom[7]      = 32'b00000000010000000110000110010011;
                     rom[8]      = 32'b00000000001100001100001001100011;
                     rom[9]      = 32'b00000010011000000000000001101111;
                     rom[10]     = 32'b01000000000100011000001000110011;
                     rom[11]     = 32'b00000000010000010100001001100011;
                     rom[12]     = 32'b00000001101000000000000001101111;
                     rom[13]     = 32'b00000000000000010011001010000011;
                     rom[14]     = 32'b00000000000100010011001100000011;
                     rom[15]     = 32'b00000000010100110100001001100011;
                     rom[16]     = 32'b00000000111000000000000001101111;
                     rom[17]     = 32'b00000000000000101000001110010011;
                     rom[18]     = 32'b00000000000000110000001010010011;
                     rom[19]     = 32'b00000000000000111000001100010011;
                     rom[20]     = 32'b00000000010100010011000000100011;
                     rom[21]     = 32'b00000000011000010011000010100011;
                     rom[22]     = 32'b00000000001000000000000001101111;
                     rom[23]     = 32'b00000000000100010000000100010011;
                     rom[24]     = 32'b11111110010111111111000001101111;
                     rom[25]     = 32'b00000000000100001000000010010011;
                     rom[26]     = 32'b00000000000000000110000100010011;
                     rom[27]     = 32'b11111101101111111111000001101111;
                     rom[28]     = 32'b00000000000000000000000000010011;
                     rom[29]     = 32'b00000000000000000011001010000011;
                     rom[30]     = 32'b00000000000100000011001100000011;
                     rom[31]     = 32'b00000000001000000011001110000011;
                     rom[32]     = 32'b00000000001100000011010000000011;
                     rom[33]     = 32'b00000000010000000011010010000011;
                     rom[34]     = 32'b00000000000000000000000000010011;
                     rom[35]     = 32'b11111111111111111111000001101111;                    
                for (i = 36; i <= 255; i=i+1) begin
                  rom[i] = 32'd0;
                end
                
      end

      always @(posedge clk) begin
          data_out <= rom[mem_address];
      end

endmodule
