module inst_memory (
  input [7:0] mem_address,
  output [31:0] data_out
);

integer i;

reg [31:0] rom [256:0];

initial  
      begin  
                  rom[0] = 32'b00000000000000000000000010000011;
                  rom[1] = 32'b00000000000000001000000100000011;
                  rom[2] = 32'b00000000000000010000000110000011;
                  rom[3] = 32'b00000000000000011000001000000011;
                  rom[4] = 32'b00000000000000100000001010000011;
                  rom[5] = 32'b00000000000000101000001100000011;
                  rom[6] = 32'b00000000000000110000001110000011;
                  rom[7] = 32'b00000000000000111000010000000011;
                  rom[8] = 32'b00000000000001000000010010000011;
                  rom[9] = 32'b00000000000001001000010100000011;
                  rom[10] = 32'b00000000000001010000010110000011;
                  rom[11] = 32'b00000000000001011000011000000011;
                  rom[12] = 32'b00000000000001100000011010000011;
                  rom[13] = 32'b00000000000001101000011100000011;
                  rom[14] = 32'b00000000000001110000011110000011;
                  rom[15] = 32'b00000000000001111000100000000011;
                  rom[16] = 32'b00000001000001111000100010110011;
                  rom[17] = 32'b00000000010001000110110000110011;
                  rom[18] = 32'b00000001000111000011000000100011;

                for (i = 19; i <= 255; i++) begin
                  rom[i] = 32'd0;
                end
                
      end

assign data_out = rom[mem_address];

endmodule
