module h3_gen (
  input  [58:0] data_i,
  input  [6:0]  seed_i,

  output [6:0]  hash_o
);

  wire [6:0] temp_hash_w;

  assign temp_hash_w = (7'd101  & {7{data_i[58]}}) ^
                       (7'd15 & {7{data_i[57]}}) ^
                       (7'd9 & {7{data_i[56]}}) ^
                       (7'd89  & {7{data_i[55]}}) ^
                       (7'd109  & {7{data_i[54]}}) ^
                       (7'd82  & {7{data_i[53]}}) ^
                       (7'd71  & {7{data_i[52]}}) ^
                       (7'd63 & {7{data_i[51]}}) ^
                       (7'd17  & {7{data_i[50]}}) ^
                       (7'd53  & {7{data_i[49]}}) ^
                       (7'd35  & {7{data_i[48]}}) ^
                       (7'd46 & {7{data_i[47]}}) ^
                       (7'd102  & {7{data_i[46]}}) ^
                       (7'd87  & {7{data_i[45]}}) ^
                       (7'd60 & {7{data_i[44]}}) ^
                       (7'd99  & {7{data_i[43]}}) ^
                       (7'd121 & {7{data_i[42]}}) ^
                       (7'd2  & {7{data_i[41]}}) ^
                       (7'd105  & {7{data_i[40]}}) ^
                       (7'd1  & {7{data_i[39]}}) ^
                       (7'd34  & {7{data_i[38]}}) ^
                       (7'd19 & {7{data_i[37]}}) ^
                       (7'd41 & {7{data_i[36]}}) ^
                       (7'd115  & {7{data_i[35]}}) ^
                       (7'd96  & {7{data_i[34]}}) ^
                       (7'd93  & {7{data_i[33]}}) ^
                       (7'd107  & {7{data_i[32]}}) ^
                       (7'd4  & {7{data_i[31]}}) ^
                       (7'd25  & {7{data_i[30]}}) ^
                       (7'd8  & {7{data_i[29]}}) ^
                       (7'd116 & {7{data_i[28]}}) ^
                       (7'd39 & {7{data_i[27]}}) ^
                       (7'd100  & {7{data_i[26]}}) ^
                       (7'd79  & {7{data_i[25]}}) ^
                       (7'd62  & {7{data_i[24]}}) ^
                       (7'd72  & {7{data_i[23]}}) ^
                       (7'd81 & {7{data_i[22]}}) ^
                       (7'd47  & {7{data_i[21]}}) ^
                       (7'd74  & {7{data_i[20]}}) ^
                       (7'd49  & {7{data_i[19]}}) ^
                       (7'd32 & {7{data_i[18]}}) ^
                       (7'd16  & {7{data_i[17]}}) ^
                       (7'd67  & {7{data_i[16]}}) ^
                       (7'd85 & {7{data_i[15]}}) ^
                       (7'd73  & {7{data_i[14]}}) ^
                       (7'd6 & {7{data_i[13]}}) ^
                       (7'd126  & {7{data_i[12]}}) ^
                       (7'd5  & {7{data_i[11]}}) ^
                       (7'd66  & {7{data_i[10]}}) ^
                       (7'd30  & {7{data_i[9]}})  ^
                       (7'd24 & {7{data_i[8]}})  ^
                       (7'd113 & {7{data_i[7]}})  ^
                       (7'd13  & {7{data_i[6]}})  ^
                       (7'd103  & {7{data_i[5]}})  ^
                       (7'd104  & {7{data_i[4]}})  ^
                       (7'd86  & {7{data_i[3]}})  ^
                       (7'd51  & {7{data_i[2]}})  ^
                       (7'd90  & {7{data_i[1]}})  ^
                       (7'd43  & {7{data_i[0]}});                

  assign hash_o = seed_i ^ temp_hash_w;
  
endmodule
