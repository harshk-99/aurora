module inst_memory (
  input clk,
  input rst,
  input [7:0] mem_address,
  input hazard,
  output reg [31:0] data_out
);

integer i;

reg [31:0] rom [256:0];

initial  
      begin  
                  rom[0]    = 32'b00000000000000000000000010000011;
                  // rom[1]    = 32'd0;
                  // rom[2]    = 32'd0;
                  // rom[3]    = 32'd0;
                  // rom[4]    = 32'd0;
                  // rom[5]    = 32'd0;
                  rom[1]    = 32'b00000000000000001000000100000011;
                  // rom[7]    = 32'd0;
                  // rom[8]    = 32'd0;
                  // rom[9]    = 32'd0;
                  // rom[10]   = 32'd0;
                  // rom[11]   = 32'd0;
                  rom[2]   = 32'b00000000000000010000000110000011;
                  // rom[13]   = 32'd0;
                  // rom[14]   = 32'd0;
                  // rom[15]   = 32'd0;
                  // rom[16]   = 32'd0;
                  // rom[17]   = 32'd0;
                  rom[3]   = 32'b00000000000000011000001000000011;
                  // rom[19]   = 32'd0;
                  // rom[20]   = 32'd0;
                  // rom[21]   = 32'd0;
                  // rom[22]   = 32'd0;
                  // rom[23]   = 32'd0;
                  rom[4]   = 32'b00000000000000100000001010000011;
                  // rom[25]   = 32'd0;
                  // rom[26]   = 32'd0;
                  // rom[27]   = 32'd0;
                  // rom[28]   = 32'd0;
                  // rom[29]   = 32'd0;
                  rom[5]   = 32'b00000000000000101000001100000011;
                  // rom[31]   = 32'd0;
                  // rom[32]   = 32'd0;
                  // rom[33]   = 32'd0;
                  // rom[34]   = 32'd0;
                  // rom[35]   = 32'd0;
                  rom[6]   = 32'b00000000000000110000001110000011;
                  // rom[37]   = 32'd0;
                  // rom[38]   = 32'd0;
                  // rom[39]   = 32'd0;
                  // rom[40]   = 32'd0;
                  // rom[41]   = 32'd0;
                  rom[7]   = 32'b00000000000000111000010000000011;
                  // rom[43]   = 32'd0;
                  // rom[44]   = 32'd0;
                  // rom[45]   = 32'd0;
                  // rom[46]   = 32'd0;
                  // rom[47]   = 32'd0;
                  rom[8]   = 32'b00000000000001000000010010000011;
                  // rom[49]   = 32'd0;
                  // rom[50]   = 32'd0;
                  // rom[51]   = 32'd0;
                  // rom[52]   = 32'd0;
                  // rom[53]   = 32'd0;
                  rom[9]   = 32'b00000000000001001000010100000011;
                  // rom[55]   = 32'd0;
                  // rom[56]   = 32'd0;
                  // rom[57]   = 32'd0;
                  // rom[58]   = 32'd0;
                  // rom[59]   = 32'd0;
                  rom[10]   = 32'b00000000000001010000010110000011;
                  // rom[61]   = 32'd0;
                  // rom[62]   = 32'd0;
                  // rom[63]   = 32'd0;
                  // rom[64]   = 32'd0;
                  // rom[65]   = 32'd0;
                  rom[11]   = 32'b00000000000001011000011000000011;
                  // rom[67]   = 32'd0;
                  // rom[68]   = 32'd0;
                  // rom[69]   = 32'd0;
                  // rom[70]   = 32'd0;
                  // rom[71]   = 32'd0;
                  rom[12]   = 32'b00000000000001100000011010000011;
                  // rom[73]   = 32'd0;
                  // rom[74]   = 32'd0;
                  // rom[75]   = 32'd0;
                  // rom[76]   = 32'd0;
                  // rom[77]   = 32'd0;
                  rom[13]   = 32'b00000000000001101000011100000011;
                  // rom[79]   = 32'd0;
                  // rom[80]   = 32'd0;
                  // rom[81]   = 32'd0;
                  // rom[82]   = 32'd0;
                  // rom[83]   = 32'd0;
                  rom[14]   = 32'b00000000000001110000011110000011;
                  // rom[85]   = 32'd0;
                  // rom[86]   = 32'd0;
                  // rom[87]   = 32'd0;
                  // rom[88]   = 32'd0;
                  // rom[89]   = 32'd0;
                  rom[15]   = 32'b00000000000001111000100000000011;
                  // rom[91]   = 32'd0;
                  // rom[92]   = 32'd0;
                  // rom[93]   = 32'd0;
                  // rom[94]   = 32'd0;
                  // rom[95]   = 32'd0;
                  rom[16]   = 32'b00000001000001111000100010110011;
                  // rom[97]   = 32'd0;
                  // rom[98]   = 32'd0;
                  // rom[99]   = 32'd0;
                  // rom[100]  = 32'd0;
                  // rom[101]  = 32'd0;
                  rom[17]  = 32'b00000000010001000110110000110011;
                  // rom[103]  = 32'd0;
                  // rom[104]  = 32'd0;
                  // rom[105]  = 32'd0;
                  // rom[106]  = 32'd0;
                  // rom[107]  = 32'd0;
                  rom[18]  = 32'b00000001000111000011000000100011;
                  // rom[109]  = 32'd0;
                  // rom[110]  = 32'd0;
                  // rom[111]  = 32'd0;
                  // rom[112]  = 32'd0;
                  // rom[113]  = 32'd0;                  
                for (i = 19; i <= 255; i=i+1) begin
                  rom[i] = 32'd0;
                end
                
      end

      always @(posedge clk) begin
        if (!rst && !hazard)
          data_out <= rom[mem_address];
        else
          data_out <= data_out;
      end

endmodule
