module inst_memory (
  input clk,
  input rst,
  input [7:0] mem_address,
  input hazard,
  output reg [31:0] data_out
);

integer i;

reg [31:0] rom [256:0];

initial  
      begin  
                  // rom[0]    = 32'b00000000000000000000000010000011;
                  // rom[1]    = 32'b00000000000000001000000100000011;
                  // rom[2]    = 32'b00000000000000010000000110000011;
                  // rom[3]    = 32'b00000000000000011000001000000011;
                  // rom[4]    = 32'b00000000000000100000001010000011;
                  // rom[5]    = 32'b00000000000000101000001100000011;      
                  // rom[6]    = 32'b00000000000000110000001110000011;                  
                  // rom[7]    = 32'b00000000000000111000010000000011;                  
                  // rom[8]    = 32'b00000000000001000000010010000011;                  
                  // rom[9]    = 32'b00000000000001001000010100000011;                  
                  // rom[10]   = 32'b00000000000001010000010110000011;                  
                  // rom[11]   = 32'b00000000000001011000011000000011;                  
                  // rom[12]   = 32'b00000000000001100000011010000011;                
                  // rom[13]   = 32'b00000000000001101000011100000011;                  
                  // rom[14]   = 32'b00000000000001110000011110000011;                  
                  // rom[15]   = 32'b00000000000001111000100000000011;                  
                  // rom[16]   = 32'b00000001000001111000100010110011;                  
                  // rom[17]   = 32'b00000000010001000110110000110011;                  
                  // rom[18]   = 32'b00000001000111000011000000100011;                  

        
                     rom[0]      = 32'b00000000000000000110010000010011;
                     rom[1]      = 32'b00000000001100000110011110010011;
                     rom[2]      = 32'b00000000111101000011000000100011;
                     rom[3]      = 32'b00000000010100000110011110010011;
                     rom[4]      = 32'b00000000111101000011000010100011;
                     rom[5]      = 32'b00000000000100000110011110010011;
                     rom[6]      = 32'b00000000111101000011000100100011;
                     rom[7]      = 32'b00000000001000000110011110010011;
                     rom[8]      = 32'b00000000111101000011000110100011;
                     rom[9]      = 32'b00000000010000000110011110010011;
                     rom[10]     = 32'b00000000111101000011001000100011;
                     rom[11]     = 32'b00000000000000000110001010010011;
                     rom[12]     = 32'b00000000000000000110001100010011;
                     rom[13]     = 32'b00000000010000000110001110010011;
                     rom[14]     = 32'b00000000011100101100001001100011;
                     rom[15]     = 32'b00000010011000000000000001101111;
                     rom[16]     = 32'b01000000010100111000111000110011;
                     rom[17]     = 32'b00000001110000110100001001100011;
                     rom[18]     = 32'b00000001101000000000000001101111;
                     rom[19]     = 32'b00000000000000110011100100000011;
                     rom[20]     = 32'b00000000000100110011100110000011;
                     rom[21]     = 32'b00000001001010011100001001100011;
                     rom[22]     = 32'b00000000111000000000000001101111;
                     rom[23]     = 32'b00000000000010010000101000010011;
                     rom[24]     = 32'b00000000000010011000100100010011;
                     rom[25]     = 32'b00000000000010100000100110010011;
                     rom[26]     = 32'b00000001001000110011000000100011;
                     rom[27]     = 32'b00000001001100110011000010100011;
                     rom[28]     = 32'b00000000001000000000000001101111;
                     rom[29]     = 32'b00000000000100110000001100010011;
                     rom[30]     = 32'b11111110010111111111000001101111;
                     rom[31]     = 32'b00000000000100101000001010010011;
                     rom[32]     = 32'b00000000000000000110001100010011;
                     rom[33]     = 32'b11111101101111111111000001101111;
                     rom[34]     = 32'b00000000000000000000000000010011;   
                for (i = 35; i <= 255; i=i+1) begin
                  rom[i] = 32'd0;
                end
                
      end

      always @(posedge clk) begin
        if (!rst && !hazard)
          data_out <= rom[mem_address];
        else
          data_out <= data_out;
      end

endmodule
